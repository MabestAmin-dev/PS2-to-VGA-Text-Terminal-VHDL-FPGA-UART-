-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type


-- entity
entity CHAR_ROM is
	port (
		clk      : in std_logic;
		addr     : in unsigned(10 downto 0);
		data     : out std_logic_vector(7 downto 0));
end CHAR_ROM;


-- architecture
architecture Behavioral of CHAR_ROM is
	type rom_t is array (0 to 2047) of std_logic_vector(7 downto 0);
	signal ROM_DATA : rom_t;

begin

	-- Read from the ROM:
	process(clk)
	begin
		if rising_edge(clk) then
			data <= ROM_DATA(to_integer(addr));
		end if;
	end process;
	
	ROM_DATA <= (
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- space
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",  -- A
		x"FF",x"00",x"00",x"FF",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",  -- B
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",  -- C
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- D
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- E
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- F
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- G
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- H
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- I
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- J
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- K
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- L
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- M
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- N
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- O
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- P
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- Q
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- R
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- S
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- T
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- U
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- V
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",  -- W
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"E0",x"E0",x"FF",x"FF",x"FF",x"E0",x"E0",x"FF",  -- X
		x"FF",x"E0",x"E0",x"FF",x"E0",x"E0",x"FF",x"FF",
		x"FF",x"FF",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",
		x"FF",x"E0",x"E0",x"FF",x"E0",x"E0",x"FF",x"FF",
		x"E0",x"E0",x"FF",x"FF",x"FF",x"E0",x"E0",x"FF",
		x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"1C",x"1C",x"FF",x"FF",x"1C",x"1C",x"FF",  -- Y
		x"FF",x"1C",x"1C",x"FF",x"FF",x"1C",x"1C",x"FF",
		x"FF",x"1C",x"1C",x"FF",x"FF",x"1C",x"1C",x"FF",
		x"FF",x"FF",x"1C",x"1C",x"1C",x"1C",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"1C",x"1C",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"1C",x"1C",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"1C",x"1C",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"FF",  -- Z
		x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"03",x"03",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",  -- Å
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",  -- Ä
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",  -- Ö
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		
		x"FF",x"FF",x"27",x"27",x"27",x"27",x"FF",x"FF",      -- PACMAN CURSOR
		x"FF",x"27",x"27",x"27",x"27",x"27",x"27",x"FF",
		x"27",x"27",x"27",x"27",x"E0",x"27",x"FF",x"FF",
		x"27",x"27",x"27",x"27",x"27",x"FF",x"FF",x"FF",
		x"27",x"27",x"27",x"27",x"27",x"FF",x"FF",x"FF",
		x"27",x"27",x"27",x"27",x"27",x"27",x"FF",x"FF",
		x"FF",x"27",x"27",x"27",x"27",x"27",x"27",x"FF",
		x"FF",x"FF",x"27",x"27",x"27",x"27",x"FF",x"FF"
	);
	
end Behavioral;

